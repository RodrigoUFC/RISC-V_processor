library verilog;
use verilog.vl_types.all;
entity Sign_Extend_tb is
end Sign_Extend_tb;
