library verilog;
use verilog.vl_types.all;
entity testbench_instruction_decoder is
end testbench_instruction_decoder;
