library verilog;
use verilog.vl_types.all;
entity mux_Branch_tb is
end mux_Branch_tb;
