library verilog;
use verilog.vl_types.all;
entity mux_ALUSrc_tb is
end mux_ALUSrc_tb;
