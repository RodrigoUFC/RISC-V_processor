library verilog;
use verilog.vl_types.all;
entity mux_MemtoReg_tb is
end mux_MemtoReg_tb;
