library verilog;
use verilog.vl_types.all;
entity mux_reg2loc_tb is
end mux_reg2loc_tb;
