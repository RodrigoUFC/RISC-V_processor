library verilog;
use verilog.vl_types.all;
entity tb_ALUControl is
end tb_ALUControl;
